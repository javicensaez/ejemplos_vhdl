library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity registro is
    Port ( entrada : in STD_LOGIC_VECTOR (15 downto 0);
           salida : out STD_LOGIC_VECTOR (15 downto 0);
           carga : in STD_LOGIC;
           clk : in STD_LOGIC;
           rst : in STD_LOGIC);
end registro;

architecture Behavioral of registro is

begin




end Behavioral;
